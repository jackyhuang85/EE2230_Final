`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:44:24 06/09/2016 
// Design Name: 
// Module Name:    music_player 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "parameters.v"
module music_player(
    input [2:0]song_sel,
    input clk_8hz,
    input rst_n,
	input pause,
	//input clk,
    output reg[19:0]note_div
    );
	reg [2:0]song;
	reg [9:0]cnt;
	reg [9:0]cnt_tmp;
	wire [2:0] song_next;
	
	always @(*) begin
		if(pause == 1'b1) note_div = 20'd0;
		else 
		case(song)
			3'd0: begin
				case (cnt)
					10'd0: 	note_div = 20'd57307;  	//4
					10'd1: 	note_div = 20'd57307;
					10'd2: 	note_div = 20'd51020;  	//5
					10'd3: 	note_div = 20'd51020;
					10'd4:	note_div = 20'd45454; 	//6
					10'd5:	note_div = 20'd45454; 
					10'd6:	note_div = 20'd57307; 	//4  
					10'd7:	note_div = 20'd57307;
					10'd8:	note_div = 20'd38168; 	//1_high
					10'd9:	note_div = 20'd38168; 
					10'd10:	note_div = 20'd38168; 
					10'd11:	note_div = 20'd38168; 
					10'd12:  note_div = 20'd45454;	//6
					10'd13:	note_div = 20'd45454;
					10'd14:	note_div = 20'd45454;
					10'd15:	note_div = 20'd45454;
					10'd16:	note_div = 20'd51020; 	//5
					10'd17:	note_div = 20'd51020; 
					10'd18:	note_div = 20'd51020; 
					10'd19:	note_div = 20'd51020; 
					10'd20:	note_div = 20'd38168; 	//1_high
					10'd21:	note_div = 20'd38168; 
					10'd22:	note_div = 20'd38168;
					10'd23:	note_div = 20'd38168;
					10'd24: 	note_div = 20'd51020; 	//5
					10'd25: 	note_div = 20'd51020; 
					10'd26: 	note_div = 20'd51020; 
					10'd27: 	note_div = 20'd51020; 
					10'd28:	note_div = 20'd57307;	//4
					10'd29:	note_div = 20'd57307;
					10'd30:	note_div = 20'd68259; 	//2
					10'd31:	note_div = 20'd68259;
					10'd32:  note_div = 20'd45454;	//6
					10'd33:	note_div = 20'd45454;
					10'd34:  note_div = 20'd45454;	
					10'd35:	note_div = 20'd45454;
					10'd36:	note_div = 20'd57307;	//4
					10'd37:	note_div = 20'd57307;
					10'd38:	note_div = 20'd57307;
					10'd39:	note_div = 20'd57307;
					10'd40:	note_div = 20'd60606;  	//3
					10'd41:	note_div = 20'd60606;
					10'd42:	note_div = 20'd60606;
					10'd43:	note_div = 20'd60606;
					10'd44:	note_div = 20'd60606;
					10'd45:	note_div = 20'd60606;
					10'd46:	note_div = 20'd60606;
					10'd47:	note_div = 20'd0;
					10'd48:	note_div = 20'd60606;	//3
					10'd48:	note_div = 20'd60606;
					10'd50:	note_div = 20'd60606;
					10'd51:	note_div = 20'd60606;
					10'd52:	note_div = 20'd68259; 	//2
					10'd53:	note_div = 20'd68259;
					10'd54:	note_div = 20'd68259; 	 
					10'd55:	note_div = 20'd68259;
					10'd56:	note_div = 20'd60606;	//3
					10'd57:	note_div = 20'd60606;
					10'd58:	note_div = 20'd60606;
					10'd59:	note_div = 20'd60606;
					10'd60:	note_div = 20'd57307;	//4
					10'd61:	note_div = 20'd57307;
					10'd62: 	note_div = 20'd51020; 	//5
					10'd63: 	note_div = 20'd51020; 
					10'd64:	note_div = 20'd76628; 	//1
					10'd65:	note_div = 20'd76628; 
					10'd66:	note_div = 20'd38168;
					10'd67:	note_div = 20'd38168;
					10'd68:	note_div = 20'd57307;	//4
					10'd69:	note_div = 20'd57307;
					10'd70:	note_div = 20'd57307;	 
					10'd71:	note_div = 20'd57307;
					10'd72: 	note_div = 20'd51020; 	//5
					10'd73: 	note_div = 20'd51020; 
					10'd74:  note_div = 20'd45454;	//6
					10'd75:	note_div = 20'd0;
					10'd76:  note_div = `A_plus4;	//6_b7
					10'd77:	note_div = 20'd45454;
					10'd78:  note_div = 20'd45454;	 
					10'd79:	note_div = 20'd45454;
					10'd80: 	note_div = 20'd40486; 	//7
					10'd81: 	note_div = 20'd40486; 
					10'd82:  note_div = 20'd45454;	//6
					10'd83:  note_div = 20'd45454;	 
					10'd84: 	note_div = 20'd51020; 	//5
					10'd85: 	note_div = 20'd51020; 
					10'd86:	note_div = 20'd57307;	//4
					10'd87:	note_div = 20'd57307;
					10'd88: 	note_div = 20'd51020; 	//5
					10'd89: 	note_div = 20'd51020; 
					10'd90: 	note_div = 20'd51020; 	 
					10'd91: 	note_div = 20'd51020; 
					10'd92: 	note_div = 20'd51020; 	 
					10'd93: 	note_div = 20'd51020; 
					10'd94: 	note_div = 20'd51020; 	 
					10'd95: 	note_div = 20'd0; 
					10'd96:	note_div = 20'd57307;	//4
					10'd97:	note_div = 20'd57307;
					10'd98: 	note_div = 20'd51020; 	//5
					10'd99: 	note_div = 20'd51020; 
					10'd100:  note_div = 20'd45454;	//6
					10'd101:  note_div = 20'd45454;	 
					10'd102:	note_div = 20'd57307;	//4
					10'd103:	note_div = 20'd57307;
					10'd104:	note_div = 20'd38168; 	//1_high
					10'd105:	note_div = 20'd38168; 	
					10'd106:	note_div = 20'd38168; 	 
					10'd107:	note_div = 20'd38168; 
					10'd108:  note_div = 20'd45454;	//6
					10'd109:  note_div = 20'd45454;	 
					10'd110:  note_div = 20'd45454;	 
					10'd111:  note_div = 20'd45454;	 
					10'd112:  note_div = 20'd45454;	 
					10'd113:  note_div = 20'd45454;	 
					10'd114:  note_div = 20'd45454;	 
					10'd115:  note_div = 20'd45454;	
					10'd116:  note_div = 20'd51020; 	//5
					10'd117:  note_div = 20'd51020; 
					10'd118:	 note_div = 20'd38168; 	//1_high
					10'd119:	 note_div = 20'd38168; 
					10'd120:  note_div = 20'd51020; 	//5
					10'd121:  note_div = 20'd51020; 
					10'd122:	note_div = 20'd57307;	//4
					10'd123:	note_div = 20'd57307;
					10'd124:	note_div = 20'd57307;	 
					10'd125:	note_div = 20'd57307;
					10'd126:	note_div = 20'd68259; 	//2
					10'd127:	note_div = 20'd68259;
					10'd128:	note_div = 20'd68259; 	 
					10'd129:	note_div = 20'd68259;
					10'd130:	note_div = 20'd60606;	//3
					10'd131:	note_div = 20'd60606;
					10'd132:	note_div = 20'd57307;	//4
					10'd133:	note_div = 20'd57307;
					10'd134:	note_div = 20'd76628; 	//1
					10'd135:	note_div = 20'd76628; 
					10'd136:	note_div = 20'd38168;
					10'd137:	note_div = 20'd38168;
					10'd138:	note_div = 20'd76628;  
					10'd139:	note_div = 20'd76628; 
					10'd140:	note_div = 20'd38168;
					10'd141:	note_div = 20'd38168;
					10'd142:	note_div = 20'd76628; 	 
					10'd143:	note_div = 20'd76628; 
					10'd144:	note_div = 20'd38168;	//1
					10'd145:	note_div = 20'd0;
					10'd146:	note_div = 20'd68259; 	//2
					10'd147:	note_div = 20'd68259;
					10'd148:	note_div = 20'd68259; 	 
					10'd149:	note_div = 20'd68259;
					10'd150:	note_div = 20'd60606;	//3
					10'd151:	note_div = 20'd60606;
					10'd152:	note_div = 20'd60606;	 
					10'd153:	note_div = 20'd60606;
					10'd154:	note_div = 20'd57307;	//4
					10'd155:	note_div = 20'd57307;
					10'd156:  note_div = 20'd51020; 	//5
					10'd157:  note_div = 20'd51020; 
					10'd158:	note_div = 20'd38168;	//1
					10'd159:	note_div = 20'd38168;	 
					10'd160:	note_div = 20'd38168;	 
					10'd161:	note_div = 20'd38168;
					10'd162:	note_div = 20'd57307;	//4
					10'd163:	note_div = 20'd57307;
					10'd164:	note_div = 20'd57307;	 
					10'd165:	note_div = 20'd57307;
					10'd166:  	note_div = 20'd51020; 	//5
					10'd167:  	note_div = 20'd51020; 
					10'd168:  	note_div = 20'd45454;	//6
					10'd169:  	note_div = 20'd45454;	 
					10'd170:  	note_div = `A_plus4;		//6_b7
					10'd171:		note_div = 20'd45454;
					10'd172:  	note_div = 20'd45454;	 
					10'd173:		note_div = 20'd45454;
					10'd174: 	note_div = 20'd40486; 	//7
					10'd175: 	note_div = 20'd40486; 
					10'd176:  	note_div = 20'd45454;	//6
					10'd177:  	note_div = 20'd45454;	 
					10'd178: 	note_div = 20'd51020; 	//5
					10'd179: 	note_div = 20'd51020; 
					10'd180:		note_div = 20'd57307;	//4
					10'd181:		note_div = 20'd57307;
					10'd182:		note_div = 20'd57307;	//4
					10'd183:		note_div = 20'd57307;
					10'd184:		note_div = 20'd57307;	 
					10'd185:		note_div = 20'd57307;
					10'd186:		note_div = 20'd57307;	 
					10'd187:		note_div = 20'd57307;
					10'd188:		note_div = 20'd57307;	 
					10'd189:		note_div = 20'd57307;
					10'd190:		note_div = 20'd57307;	 
					10'd191:		note_div = 20'd57307;
					10'd192:		note_div = 20'd57307;	 
					10'd193:		note_div = 20'd57307;
					10'd194:  	note_div = 20'd45454;	//6
					10'd195:  	note_div = 20'd45454;	 
					10'd196:  	note_div = `A_plus4;		//6_b7
					10'd197:		note_div = 20'd45454;
					10'd198:		note_div = 20'd38168; 	//1_high
					10'd199:		note_div = 20'd38168; 	
					10'd200:		note_div = 20'd38168; 	 
					10'd201:		note_div = 20'd0; 
					10'd202:		note_div = 20'd38168; 	//1_high
					10'd203:		note_div = 20'd38168; 	
					10'd204:		note_div = 20'd38168; 	 
					10'd205:		note_div = 20'd0; 
					10'd206:		note_div = 20'd38168; 	//1_high
					10'd207:		note_div = 20'd38168; 	
					10'd208:		note_div = 20'd38168; 	 
					10'd209:		note_div = 20'd0;
					10'd210:		note_div = 20'd38168; 	//1_high
					10'd211:		note_div = 20'd38168; 	
					10'd212:		note_div = 20'd38168; 	 
					10'd213:		note_div = 20'd38168; 
					10'd214:		note_div = 20'd38168; 	//1_high
					10'd215:		note_div = 20'd38168; 	
					10'd216: 	note_div = 20'd34014;	//2_high
					10'd217: 	note_div = 20'd34014;
					10'd218:		note_div = 20'd38168; 	//1_high
					10'd219:		note_div = 20'd38168; 
					10'd220:  	note_div = `A_plus4;		//6_b7
					10'd221:		note_div = 20'd0;
					10'd222:  	note_div = 20'd45454;	//6
					10'd223:  	note_div = 20'd45454;	
					10'd224:  	note_div = 20'd45454;	 
					10'd225:  	note_div = 20'd0;	
					10'd226:  	note_div = 20'd45454;	//6
					10'd227:  	note_div = 20'd45454;	
					10'd228:  	note_div = 20'd45454;	 
					10'd229:  	note_div = 20'd0;	
					10'd230:  	note_div = 20'd45454;	//6
					10'd231:  	note_div = 20'd45454;	
					10'd232:  	note_div = 20'd45454;	 
					10'd233:  	note_div = 20'd0;	
					10'd234:  	note_div = 20'd45454;	//6
					10'd235:  	note_div = 20'd0;	
					10'd236:  	note_div = `A_plus4;		//6_b7
					10'd237:		note_div = 20'd0;
					10'd238:  	note_div = 20'd45454;	//6
					10'd239:  	note_div = 20'd45454;
					10'd240: 	note_div = 20'd51020; 	//5
					10'd241: 	note_div = 20'd51020; 
					10'd242:		note_div = 20'd57307;	//4
					10'd243:		note_div = 20'd57307;
					10'd244:		note_div = 20'd60606;	//3
					10'd245:		note_div = 20'd60606;
					10'd246:		note_div = 20'd68259; 	//2
					10'd247:		note_div = 20'd68259;
					10'd248:		note_div = 20'd68259; 	 
					10'd249:		note_div = 20'd0;
					10'd250:		note_div = 20'd68259; 	//2
					10'd251:		note_div = 20'd68259;
					10'd252:		note_div = 20'd60606;	//3
					10'd253:		note_div = 20'd60606;
					10'd254:		note_div = 20'd57307;	//4
					10'd255:		note_div = 20'd57307;
					10'd256: 	note_div = 20'd51020; 	//5
					10'd257: 	note_div = 20'd51020; 
					10'd258:		note_div = 20'd38168;	//1
					10'd259:		note_div = 20'd38168;	 
					10'd260:		note_div = 20'd38168;	 
					10'd261:		note_div = 20'd38168;
					10'd262:		note_div = 20'd57307;	//4
					10'd263:		note_div = 20'd57307;
					10'd264:		note_div = 20'd57307;	 
					10'd265:		note_div = 20'd57307;
					10'd266: 	note_div = 20'd51020; 	//5
					10'd267: 	note_div = 20'd51020; 
					10'd268:  	note_div = 20'd45454;	//6
					10'd269:  	note_div = 20'd45454;
					10'd270:  	note_div = `A_plus4;		//6_b7
					10'd271:		note_div = 20'd45454;
					10'd272:  	note_div = 20'd45454;	 
					10'd273:		note_div = 20'd45454;
					10'd274: 	note_div = 20'd40486; 	//7
					10'd275: 	note_div = 20'd40486; 
					10'd276:  	note_div = 20'd45454;	//6
					10'd277:  	note_div = 20'd45454;	 
					10'd278: 	note_div = 20'd51020; 	//5
					10'd279: 	note_div = 20'd51020; 
					10'd280:		note_div = 20'd57307;	//4
					10'd281:		note_div = 20'd57307;
					10'd282: 	note_div = 20'd51020; 	//5
					10'd283: 	note_div = 20'd51020; 
					10'd284: 	note_div = 20'd51020; 	 
					10'd285: 	note_div = 20'd51020;
					10'd286: 	note_div = 20'd51020; 	 
					10'd287: 	note_div = 20'd51020; 
					10'd288: 	note_div = 20'd51020; 	 
					10'd289: 	note_div = 20'd51020;
					10'd290:		note_div = 20'd57307;	//4
					10'd291:		note_div = 20'd57307;
					10'd292: 	note_div = 20'd51020; 	//5
					10'd293: 	note_div = 20'd51020; 
					10'd294:  	note_div = 20'd45454;	//6
					10'd295:  	note_div = 20'd45454;	 
					10'd296:		note_div = 20'd57307;	//4
					10'd297:		note_div = 20'd57307;
					10'd298:		note_div = 20'd38168; 	//1_high
					10'd299:		note_div = 20'd38168; 	
					10'd300:		note_div = 20'd38168; 	 
					10'd301:		note_div = 20'd38168;
					10'd302:		note_div = 20'd38168; 	 
					10'd303:		note_div = 20'd38168;
					10'd304:  	note_div = 20'd45454;	//6
					10'd305:  	note_div = 20'd45454;	
 					10'd306: 	note_div = 20'd51020; 	//5
					10'd307: 	note_div = 20'd51020; 
					10'd308: 	note_div = 20'd51020; 	
					10'd309: 	note_div = 20'd51020; 
					10'd310:		note_div = 20'd38168; 	//1_high
					10'd311:		note_div = 20'd38168; 	
					10'd312:		note_div = 20'd38168; 	 
					10'd313:		note_div = 20'd38168;
					10'd314: 	note_div = 20'd51020; 	//5
					10'd315: 	note_div = 20'd51020; 
					10'd316: 	note_div = 20'd51020; 	
					10'd317: 	note_div = 20'd51020; 
					10'd318:		note_div = 20'd57307;	//4
					10'd319:		note_div = 20'd57307;
					10'd320:		note_div = 20'd57307;	 
					10'd321:		note_div = 20'd57307;
					10'd322:		note_div = 20'd68259; 	//2
					10'd323:		note_div = 20'd68259;
					10'd324:		note_div = 20'd68259; 	 
					10'd325:		note_div = 20'd68259;
					10'd326:		note_div = 20'd60606;	//3
					10'd327:		note_div = 20'd60606;
					10'd328:		note_div = 20'd57307;	//4
					10'd329:		note_div = 20'd57307;
					10'd330:		note_div = 20'd38168;	//1
					10'd331:		note_div = 20'd38168;	 
					10'd332:		note_div = 20'd38168;	 
					10'd333:		note_div = 20'd38168;
					10'd334:		note_div = 20'd38168;	 
					10'd335:		note_div = 20'd38168;	 
					10'd336:		note_div = 20'd38168;	 
					10'd337:		note_div = 20'd0;
					10'd338:		note_div = 20'd38168;	//1
					10'd339:		note_div = 20'd38168;	 
					10'd340:		note_div = 20'd38168;	 
					10'd341:		note_div = 20'd38168;
					10'd342:		note_div = 20'd68259; 	//2
					10'd343:		note_div = 20'd68259;
					10'd344:		note_div = 20'd68259; 	 
					10'd345:		note_div = 20'd68259;
					10'd346:		note_div = 20'd60606;	//3
					10'd347:		note_div = 20'd60606;
					10'd348:		note_div = 20'd60606;	
					10'd349:		note_div = 20'd60606;
					10'd350:		note_div = 20'd57307;	//4
					10'd351:		note_div = 20'd57307;
				   10'd352: 	note_div = 20'd51020; 	//5
					10'd353: 	note_div = 20'd51020; 
					10'd354:		note_div = 20'd38168;	//1
					10'd355:		note_div = 20'd38168;	 
					10'd356:		note_div = 20'd38168;	 
					10'd357:		note_div = 20'd38168;
					10'd358:		note_div = 20'd57307;	//4
					10'd359:		note_div = 20'd57307;
					10'd360:		note_div = 20'd57307;	 
					10'd361:		note_div = 20'd57307;
					10'd362: 	note_div = 20'd51020; 	//5
					10'd363: 	note_div = 20'd51020;
					10'd364:  	note_div = 20'd45454;	//6
					10'd365:  	note_div = 20'd45454;	
					10'd366:  	note_div = `A_plus4;		//6_b7
					10'd367:		note_div = 20'd45454;
					10'd368:  	note_div = 20'd45454;	 
					10'd369:		note_div = 20'd45454;
					10'd370: 	note_div = 20'd40486; 	//7
					10'd371: 	note_div = 20'd40486; 
					10'd372:  	note_div = 20'd45454;	//6
					10'd373:  	note_div = 20'd45454;
					10'd374: 	note_div = 20'd51020; 	//5
					10'd375: 	note_div = 20'd51020;
					10'd376:		note_div = 20'd57307;	//4
					10'd377:		note_div = 20'd57307;
					10'd378:		note_div = 20'd57307;	//4
					10'd379:		note_div = 20'd57307;
					10'd380:		note_div = 20'd57307;	 
					10'd381:		note_div = 20'd57307;
					10'd382:		note_div = 20'd57307;	 
					10'd383:		note_div = 20'd57307;
					10'd384:		note_div = 20'd57307;	 
					10'd385:		note_div = 20'd57307;
					10'd386:		note_div = 20'd57307;	 
					10'd387:		note_div = 20'd57307;
					10'd388:		note_div = 20'd57307;	 
					10'd389:		note_div = 20'd57307;
					10'd390:		note_div = 20'd57307;	
					10'd391:		note_div = 20'd57307;
					10'd392:		note_div = 20'd57307;	
					10'd393:		note_div = 20'd57307;
					10'd394:		note_div = 20'd57307;	
					10'd395:		note_div = 20'd57307;
					10'd396:		note_div = 20'd57307;	
					10'd397:		note_div = 20'd57307;
					10'd398:  	note_div = 20'd45454;	//6
					10'd399:  	note_div = 20'd45454;	 
					10'd400:  	note_div = `A_plus4;		//6_b7
					10'd401:		note_div = 20'd45454;
					10'd402:		note_div = 20'd38168; 	//1_high
					10'd403:		note_div = 20'd38168; 	
					10'd404:		note_div = 20'd38168; 	 
					10'd405:		note_div = 20'd0; 
					10'd406:		note_div = 20'd38168; 	//1_high
					10'd407:		note_div = 20'd38168; 	
					10'd408:		note_div = 20'd38168; 	 
					10'd409:		note_div = 20'd0; 
					10'd410:		note_div = 20'd38168; 	//1_high
					10'd411:		note_div = 20'd38168; 	
					10'd412:		note_div = 20'd38168; 	 
					10'd413:		note_div = 20'd0;
					10'd414:		note_div = 20'd38168; 	//1_high
					10'd415:		note_div = 20'd38168; 	
					10'd416:		note_div = 20'd38168; 	 
					10'd417:		note_div = 20'd38168; 
					10'd418:		note_div = 20'd38168; 	//1_high
					10'd419:		note_div = 20'd38168; 	
					10'd420: 	note_div = 20'd34014;	//2_high
					10'd421: 	note_div = 20'd34014;
					10'd422:		note_div = 20'd38168; 	//1_high
					10'd423:		note_div = 20'd38168; 
					10'd424:  	note_div = `A_plus4;		//6_b7
					10'd425:		note_div = 20'd0;
					10'd426:  	note_div = 20'd45454;	//6
					10'd427:  	note_div = 20'd45454;	
					10'd428:  	note_div = 20'd45454;	 
					10'd429:  	note_div = 20'd0;	
					10'd430:  	note_div = 20'd45454;	//6
					10'd431:  	note_div = 20'd45454;	
					10'd432:  	note_div = 20'd45454;	 
					10'd433:  	note_div = 20'd0;	
					10'd434:  	note_div = 20'd45454;	//6
					10'd435:  	note_div = 20'd45454;	
					10'd436:  	note_div = 20'd45454;	 
					10'd437:  	note_div = 20'd0;	
					10'd438:  	note_div = 20'd45454;	//6
					10'd439:  	note_div = 20'd0;	
					10'd440:  	note_div = `A_plus4;		//6_b7
					10'd441:		note_div = 20'd0;
					10'd442:  	note_div = 20'd45454;	//6
					10'd443:  	note_div = 20'd45454;
					10'd444: 	note_div = 20'd51020; 	//5
					10'd445: 	note_div = 20'd51020; 
					10'd446:		note_div = 20'd57307;	//4
					10'd447:		note_div = 20'd57307;
					10'd448:		note_div = 20'd60606;	//3
					10'd449:		note_div = 20'd60606;
					10'd450:		note_div = 20'd68259; 	//2
					10'd451:		note_div = 20'd68259;
					10'd452:		note_div = 20'd68259; 	 
					10'd453:		note_div = 20'd0;
					10'd454:		note_div = 20'd68259; 	//2
					10'd455:		note_div = 20'd68259;
					10'd456:		note_div = 20'd60606;	//3
					10'd457:		note_div = 20'd60606;
					10'd458:		note_div = 20'd57307;	//4
					10'd459:		note_div = 20'd57307;
					10'd460: 	note_div = 20'd51020; 	//5
					10'd461: 	note_div = 20'd51020; 
					10'd462:		note_div = 20'd38168;	//1
					10'd463:		note_div = 20'd38168;	 
					10'd464:		note_div = 20'd38168;	 
					10'd465:		note_div = 20'd38168;
					10'd466:		note_div = 20'd57307;	//4
					10'd467:		note_div = 20'd57307;
					10'd468:		note_div = 20'd57307;	 
					10'd469:		note_div = 20'd57307;
					10'd470: 	note_div = 20'd51020; 	//5
					10'd471: 	note_div = 20'd51020; 
					10'd472:  	note_div = 20'd45454;	//6
					10'd473:  	note_div = 20'd45454;
					10'd474:  	note_div = `A_plus4;		//6_b7
					10'd475:		note_div = 20'd45454;
					10'd476:  	note_div = 20'd45454;	 
					10'd477:		note_div = 20'd45454;
					10'd478: 	note_div = 20'd40486; 	//7
					10'd479: 	note_div = 20'd40486; 
					10'd480:  	note_div = 20'd45454;	//6
					10'd481:  	note_div = 20'd45454;	 
					10'd482: 	note_div = 20'd51020; 	//5
					10'd483: 	note_div = 20'd51020; 
					10'd484:		note_div = 20'd57307;	//4
					10'd485:		note_div = 20'd57307;
					10'd486: 	note_div = 20'd51020; 	//5
					10'd487: 	note_div = 20'd51020; 
					10'd488: 	note_div = 20'd51020; 	 
					10'd489: 	note_div = 20'd51020;
					10'd490: 	note_div = 20'd51020; 	 
					10'd491: 	note_div = 20'd51020; 
					10'd492: 	note_div = 20'd51020; 	 
					10'd493: 	note_div = 20'd51020;
					10'd494:		note_div = 20'd57307;	//4
					10'd495:		note_div = 20'd57307;
					10'd496: 	note_div = 20'd51020; 	//5
					10'd497: 	note_div = 20'd51020; 
					10'd498:  	note_div = 20'd45454;	//6
					10'd499:  	note_div = 20'd45454;	 
					10'd500:		note_div = 20'd57307;	//4
					10'd501:		note_div = 20'd57307;
					10'd502:		note_div = 20'd38168; 	//1_high
					10'd503:		note_div = 20'd38168; 	
					10'd504:		note_div = 20'd38168; 	 
					10'd505:		note_div = 20'd38168;
					10'd506:		note_div = 20'd38168; 	 
					10'd507:		note_div = 20'd38168;
					10'd508:  	note_div = 20'd45454;	//6
					10'd509:  	note_div = 20'd45454;	
 					10'd510: 	note_div = 20'd51020; 	//5
					10'd511: 	note_div = 20'd51020; 
					10'd512: 	note_div = 20'd51020; 	
					10'd513: 	note_div = 20'd51020; 
					10'd514:		note_div = 20'd38168; 	//1_high
					10'd515:		note_div = 20'd38168; 	
					10'd517:		note_div = 20'd38168; 	 
					10'd517:		note_div = 20'd38168;
					10'd518: 	note_div = 20'd51020; 	//5
					10'd519: 	note_div = 20'd51020; 
					10'd520: 	note_div = 20'd51020; 	
					10'd521: 	note_div = 20'd51020; 
					10'd522:		note_div = 20'd57307;	//4
					10'd523:		note_div = 20'd57307;
					10'd524:		note_div = 20'd57307;	 
					10'd525:		note_div = 20'd57307;
					10'd526:		note_div = 20'd68259; 	//2
					10'd527:		note_div = 20'd68259;
					10'd528:		note_div = 20'd68259; 	 
					10'd529:		note_div = 20'd68259;
					10'd530:		note_div = 20'd60606;	//3
					10'd531:		note_div = 20'd60606;
					10'd532:		note_div = 20'd57307;	//4
					10'd533:		note_div = 20'd57307;
					10'd534:		note_div = 20'd38168;	//1
					10'd535:		note_div = 20'd38168;	 
					10'd536:		note_div = 20'd38168;	 
					10'd537:		note_div = 20'd38168;
					10'd538:		note_div = 20'd38168;	 
					10'd539:		note_div = 20'd38168;	 
					10'd540:		note_div = 20'd38168;	 
					10'd541:		note_div = 20'd0;
					10'd542:		note_div = 20'd38168;	//1
					10'd543:		note_div = 20'd38168;	 
					10'd544:		note_div = 20'd38168;	 
					10'd545:		note_div = 20'd38168;
					10'd546:		note_div = 20'd68259; 	//2
					10'd547:		note_div = 20'd68259;
					10'd548:		note_div = 20'd68259; 	 
					10'd549:		note_div = 20'd68259;
					10'd550:		note_div = 20'd60606;	//3
					10'd551:		note_div = 20'd60606;
					10'd552:		note_div = 20'd60606;	
					10'd553:		note_div = 20'd60606;
					10'd554:		note_div = 20'd57307;	//4
					10'd555:		note_div = 20'd57307;
				   10'd556: 	note_div = 20'd51020; 	//5
					10'd557: 	note_div = 20'd51020; 
					10'd558:		note_div = 20'd38168;	//1
					10'd559:		note_div = 20'd38168;	 
					10'd560:		note_div = 20'd38168;	 
					10'd561:		note_div = 20'd38168;
					10'd562:		note_div = 20'd57307;	//4
					10'd563:		note_div = 20'd57307;
					10'd564:		note_div = 20'd57307;	 
					10'd565:		note_div = 20'd57307;
					10'd566: 	note_div = 20'd51020; 	//5
					10'd567: 	note_div = 20'd51020;
					10'd568:  	note_div = 20'd45454;	//6
					10'd569:  	note_div = 20'd45454;	
					10'd570:  	note_div = `A_plus4;		//6_b7
					10'd571:		note_div = 20'd45454;
					10'd572:  	note_div = 20'd45454;	 
					10'd573:		note_div = 20'd45454;
					10'd574: 	note_div = 20'd40486; 	//7
					10'd575: 	note_div = 20'd40486; 
					10'd576:  	note_div = 20'd45454;	//6
					10'd577:  	note_div = 20'd45454;
					10'd578: 	note_div = 20'd51020; 	//5
					10'd579: 	note_div = 20'd51020;
					10'd580:		note_div = 20'd57307;	//4
					10'd581:		note_div = 20'd57307;
					10'd582:		note_div = 20'd57307;	//4
					10'd583:		note_div = 20'd57307;
					10'd584:		note_div = 20'd57307;	 
					10'd585:		note_div = 20'd57307;
					10'd586:		note_div = 20'd57307;	 
					10'd587:		note_div = 20'd57307;
					10'd588:		note_div = 20'd57307;	 
					10'd589:		note_div = 20'd57307;
					10'd590:		note_div = 20'd57307;	 
					10'd591:		note_div = 20'd57307;
					10'd592:		note_div = 20'd57307;	 
					10'd593:		note_div = 20'd57307;
					10'd594:		note_div = 20'd57307;	
					10'd595:		note_div = 20'd57307;
					10'd596:		note_div = 20'd57307;	
					10'd597:		note_div = 20'd57307;
					10'd598:		note_div = 20'd57307;	
					10'd599:		note_div = 20'd57307;
					10'd600:		note_div = 20'd57307;	
					10'd601:		note_div = 20'd57307;
					default:		note_div = 20'd0;
				endcase
			end
		
			3'd1: begin
				case (cnt)				
					10'd0:	note_div = `E4;	//3
					10'd1:	note_div = `E4;	
					10'd2:	note_div = `D4;	//2
					10'd3:	note_div = `D4;	  
					10'd4:	note_div = `F4;	//4
					10'd5:	note_div = `F4;	 					
					10'd6:	note_div = `E4;	//3
					10'd7:	note_div = `E4;	 
					10'd8:	note_div = `E4;	//3
					10'd9:	note_div = `E4;	 
					10'd10:	note_div = `C4;	//1
					10'd11:	note_div = `C4; 					
					10'd12:	note_div = `G4;	//5
					10'd13:	note_div = `G4;	 
					10'd14:	note_div = `B4;	//7
					10'd15:	note_div = `B4;	 
					10'd16:	note_div = `C5;	//high 1
					10'd17:	note_div = `C5;
					10'd18:	note_div = `B4;	//7
					10'd19:	note_div = `B4;
					10'd20:	note_div = `G4;	//5
					10'd21:	note_div = `C4;	//1
					10'd22:	note_div = `C4;
					10'd23:	note_div = `C4;	//1
					10'd24:	note_div = 20'd0;	//1
					10'd25:	note_div = `C4;
					10'd26:	note_div = `C4;	//1
					10'd27:	note_div = 20'd0;	
					10'd28:	note_div = `C4;	//1
					10'd29:	note_div = `C4;	
					10'd30:	note_div = `A4;	//6
					10'd31:	note_div = `A4;	
					10'd32:	note_div = `A4;	//6
					10'd33:	note_div = `A4;
					10'd34:	note_div = 20'd0;	//0
					10'd35:	note_div = 20'd0;	
					10'd36:	note_div = `A4;	//6
					10'd37:	note_div = `A4;
					10'd38:	note_div = `G4;	//5
					10'd39:	note_div = 20'd0;
					10'd40:	note_div = `G4;	//5
					10'd41:	note_div = `G4;
					10'd42:	note_div = `G4;	//5
					10'd43:	note_div = 20'd0;
					10'd44:	note_div = `G4;	//5
					10'd45:	note_div = `G4;
					10'd46:	note_div = `F4;	//4
					10'd47:	note_div = `F4;	 					
					10'd48:	note_div = `E4;	//3
					10'd49:	note_div = `E4;	 
					10'd50:	note_div = `D4;	//2
					10'd51:	note_div = `D4;	  
					10'd52:	note_div = `E4;	//3
					10'd53:	note_div = `E4;	 
					10'd54:	note_div = `F4;	//4
					10'd55:	note_div = `F4;	 					
					10'd56:	note_div = `E4;	//3
					10'd57:	note_div = `E4;
					10'd58:	note_div = `E4;	//3
					10'd59:	note_div = `E4;
					10'd60:	note_div = `E4;	//3
					10'd61:	note_div = `E4;
					10'd62:	note_div = `E4;	 
					10'd63:	note_div = 20'd0;
					10'd64:	note_div = `E4;	//3
					10'd65:	note_div = `E4;
					10'd66:	note_div = `F_plus4 ;	//#4
					10'd67:	note_div = `F_plus4 ;
					10'd68:	note_div = `G_plus4 ;	//#5
					10'd69:	note_div = `G_plus4 ;
					10'd70:	note_div = `E4;	//3
					10'd71:	note_div = `E4;	 
					10'd72:	note_div = `E4;	//3
					10'd73:	note_div = `E4;
					10'd74:	note_div = `F4;	//4
					10'd75:	note_div = `F4;	
					10'd76:	note_div = `G4;	//5
					10'd77:	note_div = `G4;
					10'd78:	note_div = `B4;	//7
					10'd79:	note_div = `B4;
					10'd80:	note_div = `D5;	//high 2
					10'd81:	note_div = `D5;
					10'd82:	note_div = `B4;	//7
					10'd83:	note_div = `B4;
					10'd84:	note_div = `C5;	//high 1
					10'd85:	note_div = `C5;
					10'd86:	note_div = 20'd0;	//high 1
					10'd87:	note_div = `C5;
					10'd88:	note_div = `C5;	//high 1
					10'd89:	note_div = `C5;
					10'd90:	note_div = 20'd0;	//0
					10'd91:	note_div = 20'd0;
					10'd92:	note_div = `C5;	//high 1
					10'd93:	note_div = `C5;
					10'd94:	note_div = `C5;	//high 1
					10'd95:	note_div = `C5;
					10'd96:	note_div = `G4;	//5
					10'd97:	note_div = `G4;
					10'd98:	note_div = `G4;	//5
					10'd99:	note_div = `G4;
					10'd100:	note_div = `A4;	//6
					10'd101:	note_div = `A4;
					10'd102:	note_div = `G4;	//5
					10'd103:	note_div = `F4;	//4
					10'd104:	note_div = 20'd0;	//4
					10'd105:	note_div = `F4;
					10'd106:	note_div = `D4;	//2
					10'd107:	note_div = `D4;	  
					10'd108:	note_div = `E4;	//3
					10'd109:	note_div = `E4;	 
					10'd110:	note_div = `F4;	//4
					10'd111:	note_div = `F4;	
					10'd112:	note_div = `G4;	//5
					10'd113:	note_div = `G4;
					10'd114:	note_div = `A4;	//6
					10'd115:	note_div = `A4;	
					10'd116:	note_div = `C4;	//1
					10'd117:	note_div = `C4;
					10'd118:	note_div = `A4;	//6
					10'd119:	note_div = `A4;
					10'd120:	note_div = `A4;	 
					10'd121:	note_div = `B4;	//7
					10'd122:	note_div = 20'd0;	//7
					10'd123:	note_div = `B4;
					10'd124:	note_div = `B4;	
					10'd125:	note_div = `B4;		
					10'd126:	note_div = `E4;	//3
					10'd127:	note_div = `E4;	
					10'd128:	note_div = `D4;	//2
					10'd129:	note_div = `D4;	  
					10'd130:	note_div = `F4;	//4
					10'd131:	note_div = `F4;	 					
					10'd132:	note_div = `E4;	//3
					10'd133:	note_div = `E4;	 
					10'd134:	note_div = `E4;	//3
					10'd135:	note_div = `E4;	 
					10'd136:	note_div = `C4;	//1
					10'd137:	note_div = `C4; 					
					10'd138:	note_div = `G4;	//5
					10'd139:	note_div = `G4;	 
					10'd140:	note_div = `B4;	//7
					10'd141:	note_div = `B4;	 
					10'd142:	note_div = `C5;	//high 1
					10'd143:	note_div = `C5;
					10'd144:	note_div = `B4;	//7
					10'd145:	note_div = `B4;
					10'd146:	note_div = `G4;	//5
					10'd147:	note_div = `C4;	//1
					10'd148:	note_div = `C4;
					10'd149:	note_div = `C4;	//1
					10'd150:	note_div = 20'd0;	//1
					10'd151:	note_div = `C4;
					10'd152:	note_div = `C4;	//1
					10'd153:	note_div = 20'd0;	
					10'd154:	note_div = `C4;	//1
					10'd155:	note_div = `C4;	
					10'd156:	note_div = `A4;	//6
					10'd157:	note_div = `A4;	
					10'd158:	note_div = `A4;	//6
					10'd159:	note_div = `A4;
					10'd160:	note_div = 20'd0;	//0
					10'd161:	note_div = 20'd0;	
					10'd162:	note_div = `A4;	//6
					10'd163:	note_div = `A4;
					10'd164:	note_div = `G4;	//5
					10'd165:	note_div = 20'd0;
					10'd166:	note_div = `G4;	//5
					10'd167:	note_div = `G4;
					10'd168:	note_div = `G4;	//5
					10'd169:	note_div = 20'd0;
					10'd170:	note_div = `G4;	//5
					10'd171:	note_div = `G4;
					10'd172:	note_div = `F4;	//4
					10'd173:	note_div = `F4;	 					
					10'd174:	note_div = `E4;	//3
					10'd175:	note_div = `E4;	 
					10'd176:	note_div = `D4;	//2
					10'd177:	note_div = `D4;	  
					10'd178:	note_div = `E4;	//3
					10'd179:	note_div = `E4;	 
					10'd180:	note_div = `F4;	//4
					10'd181:	note_div = `F4;	 					
					10'd182:	note_div = `E4;	//3
					10'd183:	note_div = `E4;
					10'd184:	note_div = `E4;	//3
					10'd185:	note_div = `E4;
					10'd186:	note_div = `E4;	//3
					10'd187:	note_div = `E4;
					10'd188:	note_div = `E4;	 
					10'd189:	note_div = 20'd0;
					10'd190:	note_div = `E4;	//3
					10'd191:	note_div = `E4;
					10'd192:	note_div = `F_plus4 ;	//#4
					10'd193:	note_div = `F_plus4 ;
					10'd194:	note_div = `G_plus4 ;	//#5
					10'd195:	note_div = `G_plus4 ;
					10'd196:	note_div = `E4;	//3
					10'd197:	note_div = `E4;	 
					10'd198:	note_div = `E4;	//3
					10'd199:	note_div = `E4;
					10'd200:	note_div = `F4;	//4
					10'd201:	note_div = `F4;	
					10'd202:	note_div = `G4;	//5
					10'd203:	note_div = `G4;
					10'd204:	note_div = `B4;	//7
					10'd205:	note_div = `B4;
					10'd206:	note_div = `D5;	//high 2
					10'd207:	note_div = `D5;
					10'd208:	note_div = `B4;	//7
					10'd209:	note_div = `B4;
					10'd210:	note_div = `C5;	//high 1
					10'd211:	note_div = `C5;
					10'd212:	note_div = 20'd0;	//high 1
					10'd213:	note_div = `C5;
					10'd214:	note_div = `C5;	//high 1
					10'd215:	note_div = `C5;
					10'd216:	note_div = 20'd0;	//0
					10'd217:	note_div = 20'd0;
					10'd218:	note_div = `C5;	//high 1
					10'd219:	note_div = `C5;
					10'd220:	note_div = `C5;	//high 1
					10'd221:	note_div = `C5;
					10'd222:	note_div = `G4;	//5
					10'd223:	note_div = `G4;
					10'd224:	note_div = `G4;	//5
					10'd225:	note_div = `G4;
					10'd226:	note_div = `A4;	//6
					10'd227:	note_div = `A4;
					10'd228:	note_div = `G4;	//5
					10'd229:	note_div = `F4;	//4
					10'd230:	note_div = `F4;
					10'd231:	note_div = `A3;	//low 6
					10'd232:	note_div = `A3;
					10'd233:	note_div = `B3;	//low 7
					10'd234:	note_div = `B3;
					10'd235:	note_div = `C4;	//1
					10'd236:	note_div = `C4;	
					10'd237:	note_div = `D4;	//2
					10'd238:	note_div = `D4;	  
					10'd239:	note_div = `E4;	//3
					10'd240:	note_div = `E4;
					10'd241:	note_div = `D4;	//2
					10'd242:	note_div = `D4;
					10'd243:	note_div = `D4;	//2
					10'd244:	note_div = `D4;
					10'd245:	note_div = `D4;	 
					10'd246:	note_div = `D4;
					10'd247:	note_div = `E4;	//3
					10'd248:	note_div = `E4;
					10'd249:	note_div = `C4;	//1
					10'd250:	note_div = `C4;	
					10'd251:	note_div = `C4;	//1
					10'd252:	note_div = `C4;
					10'd253:	note_div = `C4;	 
					10'd254:	note_div = `C4;	
					default:	note_div = 20'd0;
				endcase
			end
			
			3'd2: begin
				case (cnt)
				 
					10'd0:	note_div = 20'd0;
					10'd1:	note_div = `G3;
					10'd2:	note_div = `G3;
					10'd3:	note_div = `C4;
					10'd4:	note_div = `C4;
					10'd5:	note_div = `D4;
					10'd6:	note_div = `D4;
					10'd7:	note_div = `E4;
					10'd8:	note_div = `E4;
					10'd9:	note_div = 20'd0;
					10'd10:	note_div = `E4;
					10'd11:	note_div = `E4;
					10'd12:	note_div = 20'd0;
					10'd13:	note_div = `E4;
					10'd14:	note_div = `E4;
					10'd15:	note_div = `F4;
					10'd16:	note_div = `F4;
					10'd17:	note_div = `E4;
					10'd18:	note_div = `E4;
					10'd19:	note_div = `D4;
					10'd20:	note_div = `B3;
					10'd21:	note_div = 20'd0;
					10'd22:	note_div = `B3;
					10'd23:	note_div = `D4;
					10'd24:	note_div = `D4;
					10'd25:	note_div = `C4;
					10'd26:	note_div = 20'd0;
					10'd27:	note_div = `C4;
					10'd28:	note_div = `C4;
					10'd29:	note_div = `C4;
					10'd30:	note_div = `C4;
					10'd31:	note_div = 20'd0;
					10'd32:	note_div = 20'd0;
					10'd33:	note_div = `C4;
					10'd34:	note_div = `C4;
					10'd35:	note_div = `E4;
					10'd36:	note_div = `E4;
					10'd37:	note_div = `G4;
					10'd38:	note_div = `G4;
					10'd39:	note_div = `A4;
					10'd40:	note_div = `A4;
					10'd41:	note_div = 20'd0;
					10'd42:	note_div = `A4;
					10'd43:	note_div = `A4;
					10'd44:	note_div = 20'd0;
					10'd45:	note_div = `A4;
					10'd46:	note_div = `A4;
					10'd47:	note_div = `G4;
					10'd48:	note_div = `G4;
					10'd49:	note_div = `D4;
					10'd50:	note_div = `D4;
					10'd51:	note_div = `E4;
					10'd52:	note_div = `E4;
					10'd53:	note_div = `F4;
					10'd54:	note_div = 20'd0;
					10'd55:	note_div = `F4;
					10'd56:	note_div = `E4;
					10'd57:	note_div = 20'd0;
					10'd58:	note_div = `E4;
					10'd59:	note_div = `E4;
					10'd60:	note_div = `E4;
					10'd61:	note_div = `E4;
					10'd62:	note_div = `E4;
					10'd63:	note_div = 20'd0;
					10'd64:	note_div = 20'd0;
					10'd65:	note_div = `C4;
					10'd66:	note_div = `C4;
					10'd67:	note_div = `E4;
					10'd68:	note_div = `E4;
					10'd69:	note_div = `G4;
					10'd70:	note_div = `G4;
					10'd71:	note_div = `A4;
					10'd72:	note_div = `A4;
					10'd73:	note_div = 20'd0;
					10'd74:	note_div = `A4;
					10'd75:	note_div = `A4;
					10'd76:	note_div = `A4;
					10'd77:	note_div = `A4;
					10'd78:	note_div = `A4;
					10'd79:	note_div = `B4;
					10'd80:	note_div = `B4;
					10'd81:	note_div = `A4;
					10'd82:	note_div = `A4;
					10'd83:	note_div = `G4;
					10'd84:	note_div = `F4;
					10'd85:	note_div = 20'd0;
					10'd86:	note_div = `F4;
					10'd87:	note_div = `E4;
					10'd88:	note_div = `E4;
					10'd89:	note_div = `E4;
					10'd90:	note_div = `E4;
					10'd91:	note_div = `G4;
					10'd92:	note_div = `A4;
					10'd93:	note_div = `A4;
					10'd94:	note_div = `A4;
					10'd95:	note_div = `C4;
					10'd96:	note_div = `C4;
					10'd97:	note_div = `C4;
					10'd98:	note_div = `C4;
					10'd99:	note_div = `D4;
					10'd100:	note_div = `D4;
					10'd101:	note_div = `E4;
					10'd102:	note_div = `E4;
					10'd103:	note_div = `F4;
					10'd104:	note_div = `F4;
					10'd105:	note_div = `F4;
					10'd106:	note_div = `F4;
					10'd107:	note_div = 20'd0;
					10'd108:	note_div = 20'd0;
					10'd109:	note_div = `E4;
					10'd110:	note_div = `F4;
					10'd111:	note_div = `E4;
					10'd112:	note_div = `D4;
					10'd113:	note_div = `C4;
					10'd114:	note_div = `C4;
					10'd115:	note_div = `B3;
					10'd116:	note_div = `B3;
					10'd117:	note_div = `D4;
					10'd118:	note_div = `D4;
					10'd119:	note_div = `C4;
					10'd120:	note_div = 20'd0;
					10'd121:	note_div = `C4;
					10'd122:	note_div = `C4;
					10'd123:	note_div = `C4;
					10'd124:	note_div = `C4;
					10'd125:	note_div = `C4;
					10'd126:	note_div = `C4;
					10'd127:	note_div = `C4;
					10'd128:	note_div = `C4;
				   default: note_div = 20'd0;
				endcase
			end
			
			3'd3: begin
				case (cnt)
			 
					10'd0:	note_div = `G4;
					10'd1:	note_div = `G4;
					10'd2:	note_div = `G4;
					10'd3:	note_div = `G4;
					10'd4:	note_div = `E4;
					10'd5:	note_div = `E4;
					10'd6:	note_div = `A4;
					10'd7:	note_div = `A4;
					10'd8:	note_div = `A4;
					10'd9:	note_div = `A4;
					10'd10:	note_div = `G4;
					10'd11:	note_div = `G4;
					10'd12:	note_div = `G4;
					10'd13:	note_div = `G4;
					10'd14:	note_div = `C4;
					10'd15:	note_div = `C4;
					10'd16:	note_div = `C4;
					10'd17:	note_div = `C4;
					10'd18:	note_div = `D4;
					10'd19:	note_div = `D4;
					10'd20:	note_div = `E4;
					10'd21:	note_div = `E4;
					10'd22:	note_div = `E4;
					10'd23:	note_div = `E4;
					10'd24:	note_div = `C4;
					10'd25:	note_div = `C4;
					10'd26:	note_div = `C4;
					10'd27:	note_div = `C4;
					10'd28:	note_div = `C4;
					10'd29:	note_div = `C4;
					10'd30:	note_div = `C5;
					10'd31:	note_div = `C5;
					10'd32:	note_div = `C5;
					10'd33:	note_div = `C5;
					10'd34:	note_div = `D5;
					10'd35:	note_div = `D5;
					10'd36:	note_div = `C5;
					10'd37:	note_div = `C5;
					10'd38:	note_div = `A4;
					10'd39:	note_div = `A4;
					10'd40:	note_div = `A4;
					10'd41:	note_div = `A4;
					10'd42:	note_div = `E4;
					10'd43:	note_div = `E4;
					10'd44:	note_div = `E4;
					10'd45:	note_div = `E4;
					10'd46:	note_div = `G4;
					10'd47:	note_div = `G4;
					10'd48:	note_div = `G4;
					10'd49:	note_div = `G4;
					10'd50:	note_div = `G4;
					10'd51:	note_div = `G4;
					10'd52:	note_div = `G4;
					10'd53:	note_div = `G4;
					10'd54:	note_div = `G4;
					10'd55:	note_div = `G4;
					10'd56:	note_div = `G4;
					10'd57:	note_div = `G4;
					10'd58:	note_div = `G4;
					10'd59:	note_div = `G4;
					10'd60:	note_div = `G4;
					10'd61:	note_div = `G4;
					10'd62:	note_div = `A4;
					10'd63:	note_div = `A4;
					10'd64:	note_div = `A4;
					10'd65:	note_div = `A4;
					10'd66:	note_div = `G4;
					10'd67:	note_div = `G4;
					10'd68:	note_div = `A4;
					10'd69:	note_div = `A4;
					10'd70:	note_div = `C5;
					10'd71:	note_div = `C5;
					10'd72:	note_div = `C5;
					10'd73:	note_div = `C5;
					10'd74:	note_div = `C5;
					10'd75:	note_div = `C5;
					10'd76:	note_div = `A4;
					10'd77:	note_div = `A4;
					10'd78:	note_div = `G4;
					10'd79:	note_div = `G4;
					10'd80:	note_div = `G4;
					10'd81:	note_div = `G4;
					10'd82:	note_div = `G4;
					10'd83:	note_div = `G4;
					10'd84:	note_div = `E4;
					10'd85:	note_div = `E4;
					10'd86:	note_div = `E4;
					10'd87:	note_div = `E4;
					10'd88:	note_div = `E4;
					10'd89:	note_div = `E4;
					10'd90:	note_div = `E4;
					10'd91:	note_div = 20'd0;
					10'd92:	note_div = `E4;
					10'd93:	note_div = `E4;
					10'd94:	note_div = `D4;
					10'd95:	note_div = `D4;
					10'd96:	note_div = `E4;
					10'd97:	note_div = `E4;
					10'd98:	note_div = `G4;
					10'd99:	note_div = `G4; 
					10'd100:	note_div = `E4;
					10'd101:	note_div = `E4;
					10'd102:	note_div = `E4;
					10'd103:	note_div = `E4;
					10'd104:	note_div = `D4;
					10'd105:	note_div = `D4;
					10'd106:	note_div = `D4;
					10'd107:	note_div = `D4;
					10'd108:	note_div = `C4;
					10'd109:	note_div = `C4;
					10'd110:	note_div = `C4;
					10'd111:	note_div = `C4;
					10'd112:	note_div = `E4;
					10'd113:	note_div = `E4;
					10'd114:	note_div = `E4;
					10'd115:	note_div = `E4;
					10'd116:	note_div = `D4;
					10'd117:	note_div = `D4;
					10'd118:	note_div = `D4;
					10'd119:	note_div = `D4;
					10'd120:	note_div = `D4;
					10'd121:	note_div = `D4;
					10'd122:	note_div = `D4;
					10'd123:	note_div = `D4;
					10'd124:	note_div = `D4;
					10'd125:	note_div = `D4;
					10'd126:	note_div = `D4;
					10'd127:	note_div = `D4;
					10'd128:	note_div = `D4;
					10'd129:	note_div = `D4;
					10'd130:	note_div = `G4;
					10'd131:	note_div = `G4;
					10'd132:	note_div = `G4;
					10'd133:	note_div = `G4;
					10'd134:	note_div = `E4;
					10'd135:	note_div = `E4;
					10'd136:	note_div = `A4;
					10'd137:	note_div = `A4;
					10'd138:	note_div = `A4;
					10'd139:	note_div = `A4;
					10'd140:	note_div = `G4;
					10'd141:	note_div = `G4;
					10'd142:	note_div = `G4;
					10'd143:	note_div = `G4;
					10'd144:	note_div = `C4;
					10'd145:	note_div = `C4;
					10'd146:	note_div = `C4;
					10'd147:	note_div = `C4;
					10'd148:	note_div = `D4;
					10'd149:	note_div = `D4;
					10'd150:	note_div = `E4;
					10'd151:	note_div = `E4;
					10'd152:	note_div = `E4;
					10'd153:	note_div = `E4;
					10'd154:	note_div = `C4;
					10'd155:	note_div = `C4;
					10'd156:	note_div = `C4;
					10'd157:	note_div = `C4;
					10'd158:	note_div = `C4;
					10'd159:	note_div = `C4;
					10'd160:	note_div = `C5;
					10'd170:	note_div = `C5;
					10'd171:	note_div = `C5;
					10'd172:	note_div = `C5;
					10'd173:	note_div = `D5;
					10'd174:	note_div = `D5;
					10'd175:	note_div = `C5;
					10'd176:	note_div = `C5;
					10'd177:	note_div = `A4;
					10'd178:	note_div = `A4;
					10'd179:	note_div = `A4;
					10'd180:	note_div = `A4;
					10'd181:	note_div = `E4;
					10'd182:	note_div = `E4;
					10'd183:	note_div = `E4;
					10'd184:	note_div = `E4;
					10'd185:	note_div = `G4;
					10'd186:	note_div = `G4;
					10'd187:	note_div = `G4;
					10'd188:	note_div = `G4;
					10'd189:	note_div = `G4;
					10'd190:	note_div = `G4;
					10'd191:	note_div = `G4;
					10'd192:	note_div = `G4;
					10'd193:	note_div = `G4;
					10'd194:	note_div = `G4;
					10'd195:	note_div = `G4;
					10'd196:	note_div = `G4;
					10'd197:	note_div = `G4;
					10'd198:	note_div = `G4;
					10'd199:	note_div = `G4;
					10'd200:	note_div = `G4;
					10'd201:	note_div = `A4;
					10'd202:	note_div = `A4;
					10'd203:	note_div = `A4;
					10'd204:	note_div = `A4;
					10'd205:	note_div = `G4;
					10'd206:	note_div = `G4;
					10'd207:	note_div = `A4;
					10'd208:	note_div = `A4;
					10'd209:	note_div = `C5;
					10'd210:	note_div = `C5;
					10'd211:	note_div = `C5;
					10'd212:	note_div = `C5;
					10'd213:	note_div = `C5;
					10'd214:	note_div = `C5;
					10'd215:	note_div = `A4;
					10'd216:	note_div = `A4;
					10'd217:	note_div = `G4;
					10'd218:	note_div = `G4;
					10'd219:	note_div = `G4;
					10'd220:	note_div = `G4;
					10'd221:	note_div = `G4;
					10'd222:	note_div = `G4;
					10'd223:	note_div = `E4;
					10'd224:	note_div = `E4;
					10'd225:	note_div = `E4;
					10'd226:	note_div = `E4;
					10'd227:	note_div = `E4;
					10'd228:	note_div = `E4;
					10'd229:	note_div = `E4;
					10'd230:	note_div = 20'd0;
					10'd231:	note_div = `E4;
					10'd232:	note_div = `E4;
					10'd234:	note_div = `D4;
					10'd235:	note_div = `D4;
					10'd236:	note_div = `E4;
					10'd237:	note_div = `E4;
					10'd238:	note_div = `G4;
					10'd239:	note_div = `G4; 
					10'd240:	note_div = `E4;
					10'd241:	note_div = `E4;
					10'd242:	note_div = `E4;
					10'd243:	note_div = `E4;
					10'd244:	note_div = `D4;
					10'd245:	note_div = `D4;
					10'd246:	note_div = `D4;
					10'd247:	note_div = `D4;
					10'd248:	note_div = `C4;
					10'd249:	note_div = `C4;
					10'd250:	note_div = `C4;
					10'd251:	note_div = `C4;
					10'd252:	note_div = `A3;
					10'd253:	note_div = `A3;
					10'd254:	note_div = `A3;
					10'd255:	note_div = `A3;
					10'd256:	note_div = `C4;
					10'd257:	note_div = `C4;
					10'd258:	note_div = `C4;
					10'd259:	note_div = `C4;
					10'd260:	note_div = `C4;
					10'd261:	note_div = `C4;
					10'd262:	note_div = `C4;
					10'd263:	note_div = `C4;
					10'd264:	note_div = `C4;
					10'd265:	note_div = `C4;
					10'd266:	note_div = `C4;
					10'd267:	note_div = `C4;
					10'd268:	note_div = `C4;
					10'd269:	note_div = `C4;
					10'd270:	note_div = `C4;
					10'd271:	note_div = `C4;
					10'd272:	note_div = `C4;
					10'd273:	note_div = `C4;
					default: note_div = 20'd0;
				endcase
			end
			
			3'd4: begin
				case (cnt)
				 
					10'd0:	note_div = `G5;
					10'd1:	note_div = `G5;
					10'd2:	note_div = `G5;
					10'd3:	note_div = `G5;
					10'd4:	note_div = `F5;
					10'd5:	note_div = `F5;
					10'd6:	note_div = `F5;
					10'd7:	note_div = `F5;
					10'd8:	note_div = `E5;
					10'd9:	note_div = `E5;
					10'd10:	note_div = `E5;
					10'd11:	note_div = `E5;
					10'd12:	note_div = `D5;
					10'd13:	note_div = `D5;
					10'd14:	note_div = `D5;
					10'd15:	note_div = `D5;
					10'd16:	note_div = `D5;
					10'd17:	note_div = `D5;
					10'd18:	note_div = `C5;
					10'd19:	note_div = `C5;
					10'd20:	note_div = `C5;
					10'd21:	note_div = `C5;
					10'd22:	note_div = `C5;
					10'd23:	note_div = `C5;
					10'd24:	note_div = `C5;
					10'd25:	note_div = `C5;
					10'd26:	note_div = `C5;
					10'd27:	note_div = `C5;
					10'd28:	note_div = `B4;
					10'd29:	note_div = `B4;
					10'd30:	note_div = `B4;
					10'd31:	note_div = `G4;
					10'd32:	note_div = `G4;
					10'd33:	note_div = `G4;
					10'd34:	note_div = `G4;
					10'd35:	note_div = `G4;
					10'd36:	note_div = `G4;
					10'd37:	note_div = `G4;
					10'd38:	note_div = `G4;
					10'd39:	note_div = `G4;
					10'd40:	note_div = `C5;
					10'd41:	note_div = `C5;
					10'd42:	note_div = `C5;
					10'd43:	note_div = `C5;
					10'd44:	note_div = `C5;
					10'd45:	note_div = `C5;
					10'd46:	note_div = `C5;
					10'd47:	note_div = `C5;
					10'd48:	note_div = 20'd0;
					10'd49:	note_div = `C5;
					10'd50:	note_div = `C5;
					10'd51:	note_div = `C5;
					10'd52:	note_div = `C5;
					10'd53:	note_div = `C5;
					10'd54:	note_div = `C5;
					10'd55:	note_div = `C5;
					10'd56:	note_div = `E5;
					10'd57:	note_div = `E5;
					10'd58:	note_div = `E5;
					10'd59:	note_div = `E5;
					10'd60:	note_div = `E4;
					10'd61:	note_div = `E4;
					10'd62:	note_div = `E4;
					10'd63:	note_div = `E4;
					10'd64:	note_div = `F4;
					10'd65:	note_div = `F4;
					10'd66:	note_div = `F4;
					10'd67:	note_div = `F4;
					10'd68:	note_div = `G4;
					10'd69:	note_div = `G4;
					10'd70:	note_div = `G4;
					10'd71:	note_div = `G4;
					10'd72:	note_div = `A4;
					10'd73:	note_div = `A4;
					10'd74:	note_div = `A4;
					10'd75:	note_div = `A4;
					10'd76:	note_div = `A4;
					10'd77:	note_div = `A4;
					10'd78:	note_div = `F4;
					10'd79:	note_div = `F4;
					10'd80:	note_div = `F4;
					10'd81:	note_div = `F4;
					10'd82:	note_div = `F4;
					10'd83:	note_div = `F4;
					10'd84:	note_div = `F4;
					10'd85:	note_div = `F4;
					10'd86:	note_div = `F4;
					10'd87:	note_div = `F4;
					10'd88:	note_div = `A4;
					10'd89:	note_div = `A4;
					10'd90:	note_div = `A4;
					10'd91:	note_div = `C5;
					10'd92:	note_div = 20'd0;
					10'd93:	note_div = `C5;
					10'd94:	note_div = `C5;
					10'd95:	note_div = `C5;
					10'd96:	note_div = `C5;
					10'd97:	note_div = `C5;
					10'd98:	note_div = `C5;
					10'd99:	note_div = `C5;
					10'd100:note_div = 20'd0;
					10'd101:	note_div = `C5;
					10'd102:	note_div = 20'd0;
					10'd103:	note_div = `C5;
					10'd104:	note_div = `B4;
					10'd105:	note_div = `B4;
					10'd106:	note_div = `E5;
					10'd107:	note_div = `E5;
					10'd108:	note_div = `E5;
					10'd109:	note_div = `E5;
					10'd110:	note_div = `D5;
					10'd111:	note_div = `D5;
					10'd112:	note_div = `D5;
					10'd113:	note_div = `D5;
					10'd114:	note_div = `D5;
					10'd115:	note_div = `D5;
					10'd116:	note_div = `G5;
					10'd117:	note_div = `G5;
					10'd118:	note_div = `G5;
					10'd119:	note_div = `G5;
					10'd120:	note_div = `F5;
					10'd121:	note_div = `F5;
					10'd122:	note_div = `F5;
					10'd123:	note_div = `F5;
					10'd124:	note_div = `E5;
					10'd125:	note_div = `E5;
					10'd126:	note_div = `E5;
					10'd127:	note_div = `E5;
					10'd128:	note_div = `D5;
					10'd129:	note_div = `D5;
					10'd130:	note_div = `D5;
					10'd131:	note_div = `D5;
					10'd132:	note_div = `D5;
					10'd133:	note_div = `D5;
					10'd134:	note_div = `C5;
					10'd135:	note_div = `C5;
					10'd136:	note_div = `C5;
					10'd137:	note_div = `C5;
					10'd138:	note_div = `C5;
					10'd139:	note_div = `C5;
					10'd140:	note_div = `C5;
					10'd141:	note_div = `C5;
					10'd142:	note_div = `C5;
					10'd143:	note_div = `C5;
					10'd144:	note_div = `B4;
					10'd145:	note_div = `B4;
					10'd146:	note_div = `B4;
					10'd147:	note_div = `G4;
					10'd148:	note_div = `G4;
					10'd149:	note_div = `G4;
					10'd150:	note_div = `G4;
					10'd151:	note_div = `G4;
					10'd152:	note_div = `G4;
					10'd153:	note_div = `G4;
					10'd154:	note_div = `G4;
					10'd155:	note_div = `G4;
					10'd156:	note_div = `C5;
					10'd157:	note_div = `C5;
					10'd158:	note_div = `C5;
					10'd159:	note_div = `C5;
					10'd160:	note_div = `C5;
					10'd161:	note_div = `C5;
					10'd162:	note_div = `C5;
					10'd163:	note_div = `C5;
					10'd164:	note_div = 20'd0;
					10'd165:	note_div = `C5;
					10'd166:	note_div = `C5;
					10'd167:	note_div = `C5;
					10'd168:	note_div = `C5;
					10'd169:	note_div = `C5;
					10'd170:	note_div = `C5;
					10'd171:	note_div = `C5;
					10'd172:	note_div = `E5;
					10'd173:	note_div = `E5;
					10'd174:	note_div = `E5;
					10'd175:	note_div = `E5;
					10'd176:	note_div = `E4;
					10'd177:	note_div = `E4;
					10'd178:	note_div = `E4;
					10'd179:	note_div = `E4;
					10'd180:	note_div = `F4;
					10'd181:	note_div = `F4;
					10'd182:	note_div = `F4;
					10'd183:	note_div = `F4;
					10'd184:	note_div = `G4;
					10'd185:	note_div = `G4;
					10'd186:	note_div = `G4;
					10'd187:	note_div = `G4;
					10'd188:	note_div = `A4;
					10'd189:	note_div = `A4;
					10'd190:	note_div = `A4;
					10'd191:	note_div = `A4;
					10'd192:	note_div = `A4;
					10'd193:	note_div = `A4;
					10'd194:	note_div = `F4;
					10'd195:	note_div = `F4;
					10'd196:	note_div = `F4;
					10'd197:	note_div = `F4;
					10'd198:	note_div = `F4;
					10'd199:	note_div = `F4;
					10'd200:	note_div = `F4;
					10'd201:	note_div = `F4;
					10'd202:	note_div = `F4;
					10'd203:	note_div = `F4;
					10'd204:	note_div = `A4;
					10'd205:	note_div = `A4;
					10'd206:	note_div = `A4;
					10'd207:	note_div = `C5;
					10'd208:	note_div = 20'd0;
					10'd209:	note_div = `C5;
					10'd210:	note_div = `C5;
					10'd211:	note_div = `C5;
					10'd212:	note_div = `C5;
					10'd213:	note_div = `C5;
					10'd214:	note_div = `C5;
					10'd215:	note_div = `C5;
					10'd216:	note_div = 20'd0;
					10'd217:	note_div = `C5;
					10'd218:	note_div = `C5;
					10'd219:	note_div = `A4;
					10'd220:	note_div = `A4;
					10'd221:	note_div = `A4;
					10'd222:	note_div = `A4;
					10'd223:	note_div = `A4;
					10'd224:	note_div = `A4;
					10'd225:	note_div = `E5;
					10'd226:	note_div = `E5;
					10'd227:	note_div = `E5;
					10'd228:	note_div = `E5;
					10'd229:	note_div = `D5;
					10'd230:	note_div = `D5;
					10'd231:	note_div = `D5;
					10'd232:	note_div = `B4;
					10'd233:	note_div = `B4;
					10'd234:	note_div = `B4;
					10'd235:	note_div = `B4;
					10'd236:	note_div = `B4;
					10'd237:	note_div = `D5;
					10'd238:	note_div = `D5;
					10'd239:	note_div = `D5;
					10'd240:	note_div = 20'd0;
					10'd241:	note_div = `D5;
					10'd242:	note_div = `D5;
					10'd243:	note_div = `D5;
					10'd244:	note_div = `C5;
					10'd245:	note_div = 20'd0;
					10'd246:	note_div = `C5;
					10'd247:	note_div = `C5;
					10'd248:	note_div = `C5;
					10'd249:	note_div = `C5;
					10'd250:	note_div = `C5;
					10'd251:	note_div = `C5;
					10'd252:	note_div = `C5;
					default: note_div = 20'd0;
				endcase
			end
			
			3'd5:
			begin
				case (cnt)
				 
					10'd0:	note_div = `G4;
					10'd1:	note_div = `G4;
					10'd2:	note_div = 20'd0;
					10'd3:	note_div = `G4;
					10'd4:	note_div = `E4;
					10'd5:	note_div = `E4;
					10'd6:	note_div = `D4;
					10'd7:	note_div = `D4;
					10'd8:	note_div = `D4;
					10'd9:	note_div = `D4;
					10'd10:	note_div = `C4;
					10'd11:	note_div = `C4;
					10'd12:	note_div = `C4;
					10'd13:	note_div = 20'd0;
					10'd14:	note_div = `C4;
					10'd15:	note_div = `C4;
					10'd16:	note_div = `C4;
					10'd17:	note_div = 20'd0;
					10'd18:	note_div = `C4;
					10'd19:	note_div = `C4;
					10'd20:	note_div = `C4;
					10'd21:	note_div = 20'd0;
					10'd22:	note_div = `C4;
					10'd23:	note_div = `C4;
					10'd24:	note_div = `A3;
					10'd25:	note_div = `A3;
					10'd26:	note_div = `G3;
					10'd27:	note_div = `G3;
					10'd28:	note_div = `G4;
					10'd29:	note_div = `G4;
					10'd30:	note_div = `A4;
					10'd31:	note_div = `A4;
					10'd32:	note_div = `A4;
					10'd33:	note_div = 20'd0;
					10'd34:	note_div = `A4;
					10'd35:	note_div = `A4;
					10'd36:	note_div = `A4;
					10'd37:	note_div = `A4;
					10'd38:	note_div = `A4;
					10'd39:	note_div = `A4;
					10'd40:	note_div = `C4;
					10'd41:	note_div = `C4;
					10'd42:	note_div = `D4;
					10'd43:	note_div = `D4;
					10'd44:	note_div = `E4;
					10'd45:	note_div = `E4;
					10'd46:	note_div = `G4;
					10'd47:	note_div = `G4;
					10'd48:	note_div = `G4;
					10'd49:	note_div = `G4;
					10'd50:	note_div = `G4;
					10'd51:	note_div = `G4;
					10'd52:	note_div = `G4;
					10'd53:	note_div = `G4;
					10'd54:	note_div = `C4;
					10'd55:	note_div = `C4;
					10'd56:	note_div = `C4;
					10'd57:	note_div = `C4;
					10'd58:	note_div = `D4;
					10'd59:	note_div = `D4;
					10'd60:	note_div = `D4;
					10'd61:	note_div = `D4;
					10'd62:	note_div = `D4;
					10'd63:	note_div = `D4;
					10'd64:	note_div = `D4;
					10'd65:	note_div = `D4;
					10'd66:	note_div = `D4;
					10'd67:	note_div = 20'd0;
					10'd68:	note_div = `D4;
					10'd69:	note_div = `D4;
					10'd70:	note_div = `C4;
					10'd71:	note_div = `C4;
					10'd72:	note_div = `C4;
					10'd73:	note_div = `C4;
					10'd74:	note_div = `B3;
					10'd75:	note_div = `B3;
					10'd76:	note_div = 20'd0;
					10'd77:	note_div = 20'd0;
					10'd78:	note_div = 20'd0;
					10'd79:	note_div = 20'd0;
					10'd80:	note_div = `C4;
					10'd81:	note_div = `C4;
					10'd82:	note_div = 20'd0;
					10'd83:	note_div = `C4;
					10'd84:	note_div = 20'd0;
					10'd85:	note_div = `C4;
					10'd86:	note_div = 20'd0;
					10'd87:	note_div = `C4;
					10'd88:	note_div = `C4;
					10'd89:	note_div = `A3;
					10'd90:	note_div = `A3;
					10'd91:	note_div = `G3;
					10'd92:	note_div = `G3;
					10'd93:	note_div = `G4;
					10'd94:	note_div = `G4;
					10'd95:	note_div = `A4;
					10'd96:	note_div = `A4;
					10'd97:	note_div = `A4;
					10'd98:	note_div = 20'd0;
					10'd99:	note_div = `A4; 
					10'd100:	note_div = `A4;
					10'd101:	note_div = 20'd0;
					10'd102:	note_div = `A4;
					10'd103:	note_div = `C4;
					10'd104:	note_div = `C4;
					10'd105:	note_div = 20'd0;
					10'd106:	note_div = `C4;
					10'd107:	note_div = `D4;
					10'd108:	note_div = `D4;
					10'd109:	note_div = `E4;
					10'd110:	note_div = `E4;
					10'd111:	note_div = `G4;
					10'd112:	note_div = `G4;
					10'd113:	note_div = `G4;
					10'd114:	note_div = `G4;
					10'd115:	note_div = `G3;
					10'd116:	note_div = `G3;
					10'd117:	note_div = `G4;
					10'd118:	note_div = `G4;
					10'd119:	note_div = `E4;
					10'd120:	note_div = `E4;
					10'd121:	note_div = `D4;
					10'd122:	note_div = 20'd0;
					10'd123:	note_div = `D4;
					10'd124:	note_div = `D4;
					10'd125:	note_div = `D4;
					10'd126:	note_div = `D4;
					10'd127:	note_div = `D4;
					10'd128:	note_div = `D4;
					10'd129:	note_div = `D4;
					10'd130:	note_div = `D4;
					10'd131:	note_div = `D4;
					10'd132:	note_div = `D4;
					10'd133:	note_div = `E4;
					10'd134:	note_div = `E4;
					10'd135:	note_div = `D4;
					10'd136:	note_div = `D4;
					10'd137:	note_div = `D4;
					10'd138:	note_div = `D4;
					10'd139:	note_div = `C4;
					10'd140:	note_div = `C4;
					10'd141:	note_div = `C4;
					10'd142:	note_div = `C4;
					10'd143:	note_div = `C4;
					10'd144:	note_div = 20'd0;
					10'd145:	note_div = `C4;
					10'd146:	note_div = `C4;
					10'd147:	note_div = `C4;
					10'd148:	note_div = 20'd0;
					10'd149:	note_div = `C4;
					10'd150:	note_div = `C4;
					10'd151:	note_div = 20'd0;
					10'd152:	note_div = `C4;
					10'd153:	note_div = `A3;
					10'd154:	note_div = `A3;
					10'd155:	note_div = `G3;
					10'd156:	note_div = `G3;
					10'd157:	note_div = 20'd0;
					10'd158:	note_div = `G3;
					10'd159:	note_div = `A4;
					10'd160:	note_div = `A4;
					10'd170:	note_div = `A4;
					10'd171:	note_div = `A4;
					10'd172:	note_div = 20'd0;
					10'd173:	note_div = `A4;
					10'd174:	note_div = `A4;
					10'd175:	note_div = `A4;
					10'd176:	note_div = `C4;
					10'd177:	note_div = `C4;
					10'd178:	note_div = 20'd0;
					10'd179:	note_div = `C4;
					10'd180:	note_div = `D4;
					10'd181:	note_div = `D4;
					10'd182:	note_div = `E4;
					10'd183:	note_div = `E4;
					10'd184:	note_div = `G4;
					10'd185:	note_div = `G4;
					10'd186:	note_div = `G4;
					10'd187:	note_div = 20'd0;
					10'd188:	note_div = `G4;
					10'd189:	note_div = `G4;
					10'd190:	note_div = 20'd0;
					10'd191:	note_div = `G4;
					10'd192:	note_div = `C4;
					10'd193:	note_div = `C4;
					10'd194:	note_div = `C4;
					10'd195:	note_div = `C4;
					10'd196:	note_div = `D4;
					10'd197:	note_div = `D4;
					10'd198:	note_div = `D4;
					10'd199:	note_div = `D4;
					10'd200:	note_div = `D4;
					10'd201:	note_div = `D4;
					10'd202:	note_div = `D4;
					10'd203:	note_div = `D4;
					10'd204:	note_div = `D4;
					10'd205:	note_div = `D4;
					10'd206:	note_div = `D4;
					10'd207:	note_div = `D4;
					10'd208:	note_div = `D4;
					10'd209:	note_div = `D4;
					10'd210:	note_div = `D4;
					10'd211:	note_div = `D4;
					10'd212:	note_div = `D4;
					10'd213:	note_div = `D4;
					default: note_div = 20'd0;
				endcase
			end
			
			default:
				note_div = 20'd0;
			
		endcase
	end
	
	assign song_next = song_sel;
	
	always @(posedge clk_8hz or negedge rst_n)
		if(~rst_n) song <= 3'd0;
		else song <= song_next;
	
	always @*
	begin
		if(song != song_sel)
			cnt_tmp = 10'd0;
		else if(pause == 1'b1)
			cnt_tmp = cnt;
		else 
			case(song)
			3'd0:
				if(cnt >= 10'd610) cnt_tmp = 10'd0;
				else cnt_tmp = cnt + 10'd1;
			3'd1:
				if(cnt >= 10'd260) cnt_tmp = 10'd0;
				else cnt_tmp = cnt + 10'd1;
			3'd2:
				if(cnt >= 10'd140) cnt_tmp = 10'd0;
				else cnt_tmp = cnt + 10'd1;
			3'd3:
				if(cnt >= 10'd280) cnt_tmp = 10'd0;
				else cnt_tmp = cnt + 10'd1;
			3'd4:
				if(cnt >= 10'd260) cnt_tmp = 10'd0;
				else cnt_tmp = cnt + 10'd1;
			3'd5:
				if(cnt >= 10'd220) cnt_tmp = 10'd0;
				else cnt_tmp = cnt + 10'd1;
			default:
				cnt_tmp = 10'd0;
		endcase
	end
	
	always @(posedge clk_8hz or negedge rst_n)
	begin
		if (~rst_n)	cnt <= 10'd0;
		else cnt <= cnt_tmp;
	end
endmodule
